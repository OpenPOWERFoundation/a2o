//wtf nop

module IOBUF #(
)
(
   input I,
   input T,
   inout IO,
   inout O
);

endmodule

