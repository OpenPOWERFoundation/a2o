//wtf nop

module OBUFDS #(
)
(
   input I,
   inout O,
   inout OB
);

endmodule

