//wtf doesnt do nothin!

module ISERDESE2 #(
   parameter DATA_RATE,
   parameter DATA_WIDTH,
   parameter INTERFACE_TYPE,
   parameter IOBDELAY,
   parameter NUM_CE,
   parameter SERDES_MODE
)
(
   input BITSLIP,
   input CE1,
   input CLK,
   input CLKB,
   input CLKDIV,
   input DDLY,
   input RST,
   output Q1,
   output Q2,
   output Q3,
   output Q4,
   output Q5,
   output Q6,
   output Q7,
   output Q8
);


endmodule

