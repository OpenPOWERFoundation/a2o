//wtf nop

module IOBUFDS #(
)
(
   input I,
   input T,
   inout IO,
   inout IOB
);

endmodule

