//wtf doesnt do nothin!

module OSERDESE2 #(
   parameter DATA_RATE_OQ,
   parameter DATA_RATE_TQ,
   parameter DATA_WIDTH,
   parameter SERDES_MODE,
   parameter TRISTATE_WIDTH
)
(
   input CLK,
   input CLKDIV,
   input DDLY,
   input RST,
   input D1,
   input D2,
   input D3,
   input D4,
   input D5,
   input D6,
   input D7,
   input D8,
   input OCE,
   input OFB,
   input T1,
   input TCE,
   output OQ,
   output TQ
);


endmodule

